import rv32i_types::*;

module l2_cache
(
    input clk,

    /* Signals from Arbiter */
    input rv32i_word mem_address,
    input logic [255:0] mem_wdata,
    input mem_read,
    input mem_write,

    /* Signals from P-memory */
    input pmem_resp,
    input [255:0] pmem_rdata,

    /* Signals to P-memory */
    output rv32i_word pmem_address,
    output logic [255:0] pmem_wdata,
    output logic pmem_read,
    output logic pmem_write,

    /* Signals to Arbiter */
    output logic mem_resp,
    output [255:0] mem_rdata,

	output logic is_hit
    );

logic hit_0, hit_1, hit_2, hit_3;
logic valid_out_0, dirty_out_0;
logic valid_out_1, dirty_out_1;
logic valid_out_2, dirty_out_2;
logic valid_out_3, dirty_out_3;
logic [2:0] lru_out;
logic load_data_0, load_tag_0, load_valid_0, load_dirty_0;
logic load_data_1, load_tag_1, load_valid_1, load_dirty_1;
logic load_data_2, load_tag_2, load_valid_2, load_dirty_2;
logic load_data_3, load_tag_3, load_valid_3, load_dirty_3;

logic valid_in, dirty_in;
logic [2:0] lru_in;
logic [1:0] way_sel;
logic load_lru;

logic [1:0] pmem_sel;
logic data_sel;
logic load_pmem_wdata;

assign is_hit = hit_0 | hit_1 | hit_2 | hit_3;


l2_cache_control l2_cache_control
(
    .clk,
    /* Signals from CPU */
    .mem_byte_enable(4'b1111),
    .mem_read,
    .mem_write,
    /* Signals from P-memory */
    .pmem_resp,
    /* Signals to P-memory */
    .pmem_read,
    .pmem_write,
    /* Signals to CPU */
    .mem_resp,

    /* Signal from Cache Datapath */
    .hit_0, .hit_1, .hit_2, .hit_3,

    .valid_out_0, .dirty_out_0,
    .valid_out_1, .dirty_out_1,
    .valid_out_2, .dirty_out_2,
    .valid_out_3, .dirty_out_3,

    .load_lru,
    .lru_out,
    .lru_in,

    /* Signal send to Cache Datapath */
    .load_data_0, .load_tag_0, .load_valid_0, .load_dirty_0,
    .load_data_1, .load_tag_1, .load_valid_1, .load_dirty_1,
    .load_data_2, .load_tag_2, .load_valid_2, .load_dirty_2,
    .load_data_3, .load_tag_3, .load_valid_3, .load_dirty_3,

    .valid_in,
    .dirty_in,
    .way_sel,
    .pmem_sel,
    .load_pmem_wdata,
    .data_sel
    );

l2_cache_datapath l2_cache_datapath
(
    .clk,

    /* Signals from Arbiter */
    .mem_address,       // Should be taking pmem_address from arbiter
    .mem_wdata,      // Should be taking pmem_wdata from arbiter

    /* Signals from P-memory */
    .pmem_rdata,

    /* Signals from Cache Control */
    .load_data_0, .load_tag_0, .load_valid_0, .load_dirty_0,
    .load_data_1, .load_tag_1, .load_valid_1, .load_dirty_1,
    .load_data_2, .load_tag_2, .load_valid_2, .load_dirty_2,
    .load_data_3, .load_tag_3, .load_valid_3, .load_dirty_3,

    .valid_in,
    .dirty_in,
    .way_sel,

    .load_lru, .lru_in, .lru_out,

    .pmem_sel, .data_sel, .load_pmem_wdata,

    /* Signals to P-memory */
    .pmem_address,
    .pmem_wdata,

    /* Signals to Arbiter */
    .mem_rdata,

    /* Signals generated by Cache Ways */
    .hit_0, .hit_1, .hit_2, .hit_3,

    .valid_out_0, .dirty_out_0,
    .valid_out_1, .dirty_out_1,
    .valid_out_2, .dirty_out_2,
    .valid_out_3, .dirty_out_3
    );

endmodule : l2_cache
